`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:27:11 11/01/2015 
// Design Name: 
// Module Name:    Multiplier_1 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Multiplier_1 (A, B);
	input wire [3:0] A;
	output reg [3:0] B;
	
	initial begin
		RSC(A);
	end
	
endmodule
